// cineraria_core.v

// Generated using ACDS version 15.0 153

`timescale 1 ps / 1 ps
module cineraria_core (
		input  wire        core_clk,             //      core.clk
		input  wire [9:0]  dipsw_export,         //     dipsw.export
		inout  wire [31:0] gpio0_export,         //     gpio0.export
		output wire [9:0]  led_export,           //       led.export
		output wire [15:0] led7seg_0_export,     // led7seg_0.export
		output wire [15:0] led7seg_1_export,     // led7seg_1.export
		output wire [15:0] led7seg_2_export,     // led7seg_2.export
		input  wire        pcm_clk,              //       pcm.clk
		output wire        pcm_mute,             //          .mute
		output wire        pcm_aud_l,            //          .aud_l
		output wire        pcm_aud_r,            //          .aud_r
		input  wire        peri_clk,             //      peri.clk
		inout  wire        ps2_kb_CLK,           //    ps2_kb.CLK
		inout  wire        ps2_kb_DAT,           //          .DAT
		input  wire [3:0]  psw_export,           //       psw.export
		input  wire        reset_reset_n,        //     reset.reset_n
		output wire        sd_nCS,               //        sd.nCS
		output wire        sd_SCK,               //          .SCK
		output wire        sd_SDO,               //          .SDO
		input  wire        sd_SDI,               //          .SDI
		input  wire        sd_CD,                //          .CD
		input  wire        sd_WP,                //          .WP
		output wire [12:0] sdr_addr,             //       sdr.addr
		output wire [1:0]  sdr_ba,               //          .ba
		output wire        sdr_cas_n,            //          .cas_n
		output wire        sdr_cke,              //          .cke
		output wire        sdr_cs_n,             //          .cs_n
		inout  wire [15:0] sdr_dq,               //          .dq
		output wire [1:0]  sdr_dqm,              //          .dqm
		output wire        sdr_ras_n,            //          .ras_n
		output wire        sdr_we_n,             //          .we_n
		output wire        usb_test_dataouttick, //       usb.test_dataouttick
		output wire        usb_test_dataintick,  //          .test_dataintick
		input  wire        usb_usbclk_48mhz,     //          .usbclk_48mhz
		inout  wire        usb_usb_dp,           //          .usb_dp
		inout  wire        usb_usb_dm,           //          .usb_dm
		output wire        usb_usb_oe_n,         //          .usb_oe_n
		output wire        usb_usb_fullspeed,    //          .usb_fullspeed
		input  wire        vga_clk,              //       vga.clk
		output wire [4:0]  vga_rout,             //          .rout
		output wire [4:0]  vga_gout,             //          .gout
		output wire [4:0]  vga_bout,             //          .bout
		output wire        vga_hsync_n,          //          .hsync_n
		output wire        vga_vsync_n,          //          .vsync_n
		output wire        vga_enable            //          .enable
	);

	wire  [31:0] nios2_fast_custom_instruction_master_multi_dataa;                              // nios2_fast:A_ci_multi_dataa -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_dataa
	wire         nios2_fast_custom_instruction_master_multi_writerc;                            // nios2_fast:A_ci_multi_writerc -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_writerc
	wire  [31:0] nios2_fast_custom_instruction_master_multi_result;                             // nios2_fast_custom_instruction_master_translator:ci_slave_multi_result -> nios2_fast:A_ci_multi_result
	wire         nios2_fast_custom_instruction_master_clk;                                      // nios2_fast:A_ci_multi_clock -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] nios2_fast_custom_instruction_master_multi_datab;                              // nios2_fast:A_ci_multi_datab -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_datab
	wire         nios2_fast_custom_instruction_master_start;                                    // nios2_fast:A_ci_multi_start -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_start
	wire   [4:0] nios2_fast_custom_instruction_master_multi_b;                                  // nios2_fast:A_ci_multi_b -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_b
	wire   [4:0] nios2_fast_custom_instruction_master_multi_c;                                  // nios2_fast:A_ci_multi_c -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_c
	wire         nios2_fast_custom_instruction_master_reset_req;                                // nios2_fast:A_ci_multi_reset_req -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         nios2_fast_custom_instruction_master_done;                                     // nios2_fast_custom_instruction_master_translator:ci_slave_multi_done -> nios2_fast:A_ci_multi_done
	wire   [4:0] nios2_fast_custom_instruction_master_multi_a;                                  // nios2_fast:A_ci_multi_a -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_a
	wire         nios2_fast_custom_instruction_master_clk_en;                                   // nios2_fast:A_ci_multi_clk_en -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_clken
	wire         nios2_fast_custom_instruction_master_reset;                                    // nios2_fast:A_ci_multi_reset -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_reset
	wire         nios2_fast_custom_instruction_master_multi_readrb;                             // nios2_fast:A_ci_multi_readrb -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_readrb
	wire         nios2_fast_custom_instruction_master_multi_readra;                             // nios2_fast:A_ci_multi_readra -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_readra
	wire   [7:0] nios2_fast_custom_instruction_master_multi_n;                                  // nios2_fast:A_ci_multi_n -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_n
	wire         nios2_fast_custom_instruction_master_translator_multi_ci_master_readra;        // nios2_fast_custom_instruction_master_translator:multi_ci_master_readra -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] nios2_fast_custom_instruction_master_translator_multi_ci_master_a;             // nios2_fast_custom_instruction_master_translator:multi_ci_master_a -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] nios2_fast_custom_instruction_master_translator_multi_ci_master_b;             // nios2_fast_custom_instruction_master_translator:multi_ci_master_b -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         nios2_fast_custom_instruction_master_translator_multi_ci_master_clk;           // nios2_fast_custom_instruction_master_translator:multi_ci_master_clk -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios2_fast_custom_instruction_master_translator_multi_ci_master_readrb;        // nios2_fast_custom_instruction_master_translator:multi_ci_master_readrb -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] nios2_fast_custom_instruction_master_translator_multi_ci_master_c;             // nios2_fast_custom_instruction_master_translator:multi_ci_master_c -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         nios2_fast_custom_instruction_master_translator_multi_ci_master_start;         // nios2_fast_custom_instruction_master_translator:multi_ci_master_start -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         nios2_fast_custom_instruction_master_translator_multi_ci_master_reset_req;     // nios2_fast_custom_instruction_master_translator:multi_ci_master_reset_req -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios2_fast_custom_instruction_master_translator_multi_ci_master_done;          // nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_done -> nios2_fast_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios2_fast_custom_instruction_master_translator_multi_ci_master_n;             // nios2_fast_custom_instruction_master_translator:multi_ci_master_n -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] nios2_fast_custom_instruction_master_translator_multi_ci_master_result;        // nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_result -> nios2_fast_custom_instruction_master_translator:multi_ci_master_result
	wire         nios2_fast_custom_instruction_master_translator_multi_ci_master_clk_en;        // nios2_fast_custom_instruction_master_translator:multi_ci_master_clken -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] nios2_fast_custom_instruction_master_translator_multi_ci_master_datab;         // nios2_fast_custom_instruction_master_translator:multi_ci_master_datab -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] nios2_fast_custom_instruction_master_translator_multi_ci_master_dataa;         // nios2_fast_custom_instruction_master_translator:multi_ci_master_dataa -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios2_fast_custom_instruction_master_translator_multi_ci_master_reset;         // nios2_fast_custom_instruction_master_translator:multi_ci_master_reset -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         nios2_fast_custom_instruction_master_translator_multi_ci_master_writerc;       // nios2_fast_custom_instruction_master_translator:multi_ci_master_writerc -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_readra;         // nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_readra -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_a;              // nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_a -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_b;              // nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_b -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_readrb;         // nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_readrb -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_c;              // nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_c -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_clk;            // nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_clk -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_ipending;       // nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_ipending -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_start;          // nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_start -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_reset_req;      // nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_done;           // nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_done -> nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_n;              // nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_n -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_result;         // nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_result -> nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_estatus;        // nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_estatus -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_clk_en;         // nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_clken -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_datab;          // nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_datab -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_dataa;          // nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_dataa -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_reset;          // nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_reset -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_writerc;        // nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_writerc -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_result; // nios_custom_instr_floating_point_0:result -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_clk;    // nios2_fast_custom_instruction_master_multi_slave_translator0:ci_master_clk -> nios_custom_instr_floating_point_0:clk
	wire         nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_clk_en; // nios2_fast_custom_instruction_master_multi_slave_translator0:ci_master_clken -> nios_custom_instr_floating_point_0:clk_en
	wire  [31:0] nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_datab;  // nios2_fast_custom_instruction_master_multi_slave_translator0:ci_master_datab -> nios_custom_instr_floating_point_0:datab
	wire  [31:0] nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_dataa;  // nios2_fast_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> nios_custom_instr_floating_point_0:dataa
	wire         nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_start;  // nios2_fast_custom_instruction_master_multi_slave_translator0:ci_master_start -> nios_custom_instr_floating_point_0:start
	wire         nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_reset;  // nios2_fast_custom_instruction_master_multi_slave_translator0:ci_master_reset -> nios_custom_instr_floating_point_0:reset
	wire         nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_done;   // nios_custom_instr_floating_point_0:done -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire   [1:0] nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_n;      // nios2_fast_custom_instruction_master_multi_slave_translator0:ci_master_n -> nios_custom_instr_floating_point_0:n
	wire         nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_readra;         // nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_readra -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_readra
	wire   [4:0] nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_a;              // nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_a -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_a
	wire   [4:0] nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_b;              // nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_b -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_b
	wire         nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_readrb;         // nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_readrb -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_readrb
	wire   [4:0] nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_c;              // nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_c -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_c
	wire         nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_clk;            // nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_clk -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_clk
	wire  [31:0] nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_ipending;       // nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_ipending -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_ipending
	wire         nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_start;          // nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_start -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_start
	wire         nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_reset_req;      // nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_reset_req -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_reset_req
	wire         nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_done;           // nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_done -> nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_done
	wire   [7:0] nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_n;              // nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_n -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_n
	wire  [31:0] nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_result;         // nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_result -> nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_result
	wire         nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_estatus;        // nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_estatus -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_estatus
	wire         nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_clk_en;         // nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_clken -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_clken
	wire  [31:0] nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_datab;          // nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_datab -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_datab
	wire  [31:0] nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_dataa;          // nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_dataa -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_dataa
	wire         nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_reset;          // nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_reset -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_reset
	wire         nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_writerc;        // nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_writerc -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_writerc
	wire  [31:0] nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_result; // pixelsimd:result -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_master_result
	wire         nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_clk;    // nios2_fast_custom_instruction_master_multi_slave_translator1:ci_master_clk -> pixelsimd:clk
	wire         nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_clk_en; // nios2_fast_custom_instruction_master_multi_slave_translator1:ci_master_clken -> pixelsimd:clk_en
	wire  [31:0] nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_datab;  // nios2_fast_custom_instruction_master_multi_slave_translator1:ci_master_datab -> pixelsimd:datab
	wire  [31:0] nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_dataa;  // nios2_fast_custom_instruction_master_multi_slave_translator1:ci_master_dataa -> pixelsimd:dataa
	wire         nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_start;  // nios2_fast_custom_instruction_master_multi_slave_translator1:ci_master_start -> pixelsimd:start
	wire         nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_reset;  // nios2_fast_custom_instruction_master_multi_slave_translator1:ci_master_reset -> pixelsimd:reset
	wire         nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_done;   // pixelsimd:done -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_master_done
	wire   [2:0] nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_n;      // nios2_fast_custom_instruction_master_multi_slave_translator1:ci_master_n -> pixelsimd:n
	wire  [31:0] nios2_fast_data_master_readdata;                                               // mm_interconnect_0:nios2_fast_data_master_readdata -> nios2_fast:d_readdata
	wire         nios2_fast_data_master_waitrequest;                                            // mm_interconnect_0:nios2_fast_data_master_waitrequest -> nios2_fast:d_waitrequest
	wire         nios2_fast_data_master_debugaccess;                                            // nios2_fast:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_fast_data_master_debugaccess
	wire  [28:0] nios2_fast_data_master_address;                                                // nios2_fast:d_address -> mm_interconnect_0:nios2_fast_data_master_address
	wire   [3:0] nios2_fast_data_master_byteenable;                                             // nios2_fast:d_byteenable -> mm_interconnect_0:nios2_fast_data_master_byteenable
	wire         nios2_fast_data_master_read;                                                   // nios2_fast:d_read -> mm_interconnect_0:nios2_fast_data_master_read
	wire         nios2_fast_data_master_readdatavalid;                                          // mm_interconnect_0:nios2_fast_data_master_readdatavalid -> nios2_fast:d_readdatavalid
	wire         nios2_fast_data_master_write;                                                  // nios2_fast:d_write -> mm_interconnect_0:nios2_fast_data_master_write
	wire  [31:0] nios2_fast_data_master_writedata;                                              // nios2_fast:d_writedata -> mm_interconnect_0:nios2_fast_data_master_writedata
	wire   [3:0] nios2_fast_data_master_burstcount;                                             // nios2_fast:d_burstcount -> mm_interconnect_0:nios2_fast_data_master_burstcount
	wire  [31:0] nios2_fast_instruction_master_readdata;                                        // mm_interconnect_0:nios2_fast_instruction_master_readdata -> nios2_fast:i_readdata
	wire         nios2_fast_instruction_master_waitrequest;                                     // mm_interconnect_0:nios2_fast_instruction_master_waitrequest -> nios2_fast:i_waitrequest
	wire  [27:0] nios2_fast_instruction_master_address;                                         // nios2_fast:i_address -> mm_interconnect_0:nios2_fast_instruction_master_address
	wire         nios2_fast_instruction_master_read;                                            // nios2_fast:i_read -> mm_interconnect_0:nios2_fast_instruction_master_read
	wire         nios2_fast_instruction_master_readdatavalid;                                   // mm_interconnect_0:nios2_fast_instruction_master_readdatavalid -> nios2_fast:i_readdatavalid
	wire   [3:0] nios2_fast_instruction_master_burstcount;                                      // nios2_fast:i_burstcount -> mm_interconnect_0:nios2_fast_instruction_master_burstcount
	wire         vga_m1_waitrequest;                                                            // mm_interconnect_0:vga_m1_waitrequest -> vga:avm_m1_waitrequest
	wire  [31:0] vga_m1_readdata;                                                               // mm_interconnect_0:vga_m1_readdata -> vga:avm_m1_readdata
	wire  [31:0] vga_m1_address;                                                                // vga:avm_m1_address -> mm_interconnect_0:vga_m1_address
	wire         vga_m1_read;                                                                   // vga:avm_m1_read -> mm_interconnect_0:vga_m1_read
	wire         vga_m1_readdatavalid;                                                          // mm_interconnect_0:vga_m1_readdatavalid -> vga:avm_m1_readdatavalid
	wire   [9:0] vga_m1_burstcount;                                                             // vga:avm_m1_burstcount -> mm_interconnect_0:vga_m1_burstcount
	wire  [31:0] mm_interconnect_0_nios2_fast_debug_mem_slave_readdata;                         // nios2_fast:debug_mem_slave_readdata -> mm_interconnect_0:nios2_fast_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_fast_debug_mem_slave_waitrequest;                      // nios2_fast:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_fast_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_fast_debug_mem_slave_debugaccess;                      // mm_interconnect_0:nios2_fast_debug_mem_slave_debugaccess -> nios2_fast:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_fast_debug_mem_slave_address;                          // mm_interconnect_0:nios2_fast_debug_mem_slave_address -> nios2_fast:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_fast_debug_mem_slave_read;                             // mm_interconnect_0:nios2_fast_debug_mem_slave_read -> nios2_fast:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_fast_debug_mem_slave_byteenable;                       // mm_interconnect_0:nios2_fast_debug_mem_slave_byteenable -> nios2_fast:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_fast_debug_mem_slave_write;                            // mm_interconnect_0:nios2_fast_debug_mem_slave_write -> nios2_fast:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_fast_debug_mem_slave_writedata;                        // mm_interconnect_0:nios2_fast_debug_mem_slave_writedata -> nios2_fast:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_peripherals_bridge_s0_readdata;                              // peripherals_bridge:s0_readdata -> mm_interconnect_0:peripherals_bridge_s0_readdata
	wire         mm_interconnect_0_peripherals_bridge_s0_waitrequest;                           // peripherals_bridge:s0_waitrequest -> mm_interconnect_0:peripherals_bridge_s0_waitrequest
	wire         mm_interconnect_0_peripherals_bridge_s0_debugaccess;                           // mm_interconnect_0:peripherals_bridge_s0_debugaccess -> peripherals_bridge:s0_debugaccess
	wire  [23:0] mm_interconnect_0_peripherals_bridge_s0_address;                               // mm_interconnect_0:peripherals_bridge_s0_address -> peripherals_bridge:s0_address
	wire         mm_interconnect_0_peripherals_bridge_s0_read;                                  // mm_interconnect_0:peripherals_bridge_s0_read -> peripherals_bridge:s0_read
	wire   [3:0] mm_interconnect_0_peripherals_bridge_s0_byteenable;                            // mm_interconnect_0:peripherals_bridge_s0_byteenable -> peripherals_bridge:s0_byteenable
	wire         mm_interconnect_0_peripherals_bridge_s0_readdatavalid;                         // peripherals_bridge:s0_readdatavalid -> mm_interconnect_0:peripherals_bridge_s0_readdatavalid
	wire         mm_interconnect_0_peripherals_bridge_s0_write;                                 // mm_interconnect_0:peripherals_bridge_s0_write -> peripherals_bridge:s0_write
	wire  [31:0] mm_interconnect_0_peripherals_bridge_s0_writedata;                             // mm_interconnect_0:peripherals_bridge_s0_writedata -> peripherals_bridge:s0_writedata
	wire   [0:0] mm_interconnect_0_peripherals_bridge_s0_burstcount;                            // mm_interconnect_0:peripherals_bridge_s0_burstcount -> peripherals_bridge:s0_burstcount
	wire         mm_interconnect_0_sdram_s1_chipselect;                                         // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                           // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                        // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                            // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                               // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                         // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                      // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                              // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                          // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_bootmem_s1_chipselect;                                       // mm_interconnect_0:bootmem_s1_chipselect -> bootmem:chipselect
	wire  [31:0] mm_interconnect_0_bootmem_s1_readdata;                                         // bootmem:readdata -> mm_interconnect_0:bootmem_s1_readdata
	wire  [13:0] mm_interconnect_0_bootmem_s1_address;                                          // mm_interconnect_0:bootmem_s1_address -> bootmem:address
	wire   [3:0] mm_interconnect_0_bootmem_s1_byteenable;                                       // mm_interconnect_0:bootmem_s1_byteenable -> bootmem:byteenable
	wire         mm_interconnect_0_bootmem_s1_write;                                            // mm_interconnect_0:bootmem_s1_write -> bootmem:write
	wire  [31:0] mm_interconnect_0_bootmem_s1_writedata;                                        // mm_interconnect_0:bootmem_s1_writedata -> bootmem:writedata
	wire         mm_interconnect_0_bootmem_s1_clken;                                            // mm_interconnect_0:bootmem_s1_clken -> bootmem:clken
	wire         peripherals_bridge_m0_waitrequest;                                             // mm_interconnect_1:peripherals_bridge_m0_waitrequest -> peripherals_bridge:m0_waitrequest
	wire  [31:0] peripherals_bridge_m0_readdata;                                                // mm_interconnect_1:peripherals_bridge_m0_readdata -> peripherals_bridge:m0_readdata
	wire         peripherals_bridge_m0_debugaccess;                                             // peripherals_bridge:m0_debugaccess -> mm_interconnect_1:peripherals_bridge_m0_debugaccess
	wire  [23:0] peripherals_bridge_m0_address;                                                 // peripherals_bridge:m0_address -> mm_interconnect_1:peripherals_bridge_m0_address
	wire         peripherals_bridge_m0_read;                                                    // peripherals_bridge:m0_read -> mm_interconnect_1:peripherals_bridge_m0_read
	wire   [3:0] peripherals_bridge_m0_byteenable;                                              // peripherals_bridge:m0_byteenable -> mm_interconnect_1:peripherals_bridge_m0_byteenable
	wire         peripherals_bridge_m0_readdatavalid;                                           // mm_interconnect_1:peripherals_bridge_m0_readdatavalid -> peripherals_bridge:m0_readdatavalid
	wire  [31:0] peripherals_bridge_m0_writedata;                                               // peripherals_bridge:m0_writedata -> mm_interconnect_1:peripherals_bridge_m0_writedata
	wire         peripherals_bridge_m0_write;                                                   // peripherals_bridge:m0_write -> mm_interconnect_1:peripherals_bridge_m0_write
	wire   [0:0] peripherals_bridge_m0_burstcount;                                              // peripherals_bridge:m0_burstcount -> mm_interconnect_1:peripherals_bridge_m0_burstcount
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;                      // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;                        // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest;                     // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;                         // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;                            // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;                           // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;                       // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_1_ps2_kb_avalon_ps2_slave_chipselect;                          // mm_interconnect_1:ps2_kb_avalon_ps2_slave_chipselect -> ps2_kb:chipselect
	wire  [31:0] mm_interconnect_1_ps2_kb_avalon_ps2_slave_readdata;                            // ps2_kb:readdata -> mm_interconnect_1:ps2_kb_avalon_ps2_slave_readdata
	wire         mm_interconnect_1_ps2_kb_avalon_ps2_slave_waitrequest;                         // ps2_kb:waitrequest -> mm_interconnect_1:ps2_kb_avalon_ps2_slave_waitrequest
	wire   [0:0] mm_interconnect_1_ps2_kb_avalon_ps2_slave_address;                             // mm_interconnect_1:ps2_kb_avalon_ps2_slave_address -> ps2_kb:address
	wire         mm_interconnect_1_ps2_kb_avalon_ps2_slave_read;                                // mm_interconnect_1:ps2_kb_avalon_ps2_slave_read -> ps2_kb:read
	wire   [3:0] mm_interconnect_1_ps2_kb_avalon_ps2_slave_byteenable;                          // mm_interconnect_1:ps2_kb_avalon_ps2_slave_byteenable -> ps2_kb:byteenable
	wire         mm_interconnect_1_ps2_kb_avalon_ps2_slave_write;                               // mm_interconnect_1:ps2_kb_avalon_ps2_slave_write -> ps2_kb:write
	wire  [31:0] mm_interconnect_1_ps2_kb_avalon_ps2_slave_writedata;                           // mm_interconnect_1:ps2_kb_avalon_ps2_slave_writedata -> ps2_kb:writedata
	wire  [31:0] mm_interconnect_1_epcq_avl_csr_readdata;                                       // epcq:avl_csr_rddata -> mm_interconnect_1:epcq_avl_csr_readdata
	wire         mm_interconnect_1_epcq_avl_csr_waitrequest;                                    // epcq:avl_csr_waitrequest -> mm_interconnect_1:epcq_avl_csr_waitrequest
	wire   [2:0] mm_interconnect_1_epcq_avl_csr_address;                                        // mm_interconnect_1:epcq_avl_csr_address -> epcq:avl_csr_addr
	wire         mm_interconnect_1_epcq_avl_csr_read;                                           // mm_interconnect_1:epcq_avl_csr_read -> epcq:avl_csr_read
	wire         mm_interconnect_1_epcq_avl_csr_readdatavalid;                                  // epcq:avl_csr_rddata_valid -> mm_interconnect_1:epcq_avl_csr_readdatavalid
	wire         mm_interconnect_1_epcq_avl_csr_write;                                          // mm_interconnect_1:epcq_avl_csr_write -> epcq:avl_csr_write
	wire  [31:0] mm_interconnect_1_epcq_avl_csr_writedata;                                      // mm_interconnect_1:epcq_avl_csr_writedata -> epcq:avl_csr_wrdata
	wire  [31:0] mm_interconnect_1_epcq_avl_mem_readdata;                                       // epcq:avl_mem_rddata -> mm_interconnect_1:epcq_avl_mem_readdata
	wire         mm_interconnect_1_epcq_avl_mem_waitrequest;                                    // epcq:avl_mem_waitrequest -> mm_interconnect_1:epcq_avl_mem_waitrequest
	wire  [20:0] mm_interconnect_1_epcq_avl_mem_address;                                        // mm_interconnect_1:epcq_avl_mem_address -> epcq:avl_mem_addr
	wire         mm_interconnect_1_epcq_avl_mem_read;                                           // mm_interconnect_1:epcq_avl_mem_read -> epcq:avl_mem_read
	wire   [3:0] mm_interconnect_1_epcq_avl_mem_byteenable;                                     // mm_interconnect_1:epcq_avl_mem_byteenable -> epcq:avl_mem_byteenable
	wire         mm_interconnect_1_epcq_avl_mem_readdatavalid;                                  // epcq:avl_mem_rddata_valid -> mm_interconnect_1:epcq_avl_mem_readdatavalid
	wire         mm_interconnect_1_epcq_avl_mem_write;                                          // mm_interconnect_1:epcq_avl_mem_write -> epcq:avl_mem_write
	wire  [31:0] mm_interconnect_1_epcq_avl_mem_writedata;                                      // mm_interconnect_1:epcq_avl_mem_writedata -> epcq:avl_mem_wrdata
	wire   [6:0] mm_interconnect_1_epcq_avl_mem_burstcount;                                     // mm_interconnect_1:epcq_avl_mem_burstcount -> epcq:avl_mem_burstcount
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;                                // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;                                 // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_1_pcm_s0_readdata;                                             // pcm:avs_readdata -> mm_interconnect_1:pcm_s0_readdata
	wire   [1:0] mm_interconnect_1_pcm_s0_address;                                              // mm_interconnect_1:pcm_s0_address -> pcm:avs_address
	wire         mm_interconnect_1_pcm_s0_read;                                                 // mm_interconnect_1:pcm_s0_read -> pcm:avs_read
	wire         mm_interconnect_1_pcm_s0_write;                                                // mm_interconnect_1:pcm_s0_write -> pcm:avs_write
	wire  [31:0] mm_interconnect_1_pcm_s0_writedata;                                            // mm_interconnect_1:pcm_s0_writedata -> pcm:avs_writedata
	wire  [31:0] mm_interconnect_1_vga_s1_readdata;                                             // vga:avs_s1_readdata -> mm_interconnect_1:vga_s1_readdata
	wire   [1:0] mm_interconnect_1_vga_s1_address;                                              // mm_interconnect_1:vga_s1_address -> vga:avs_s1_address
	wire         mm_interconnect_1_vga_s1_read;                                                 // mm_interconnect_1:vga_s1_read -> vga:avs_s1_read
	wire         mm_interconnect_1_vga_s1_write;                                                // mm_interconnect_1:vga_s1_write -> vga:avs_s1_write
	wire  [31:0] mm_interconnect_1_vga_s1_writedata;                                            // mm_interconnect_1:vga_s1_writedata -> vga:avs_s1_writedata
	wire         mm_interconnect_1_usb_s1_chipselect;                                           // mm_interconnect_1:usb_s1_chipselect -> usb:avs_s1_chipselect
	wire   [7:0] mm_interconnect_1_usb_s1_readdata;                                             // usb:avs_s1_readdata -> mm_interconnect_1:usb_s1_readdata
	wire         mm_interconnect_1_usb_s1_waitrequest;                                          // usb:avs_s1_waitrequest -> mm_interconnect_1:usb_s1_waitrequest
	wire   [7:0] mm_interconnect_1_usb_s1_address;                                              // mm_interconnect_1:usb_s1_address -> usb:avs_s1_address
	wire         mm_interconnect_1_usb_s1_read;                                                 // mm_interconnect_1:usb_s1_read -> usb:avs_s1_read
	wire         mm_interconnect_1_usb_s1_write;                                                // mm_interconnect_1:usb_s1_write -> usb:avs_s1_write
	wire   [7:0] mm_interconnect_1_usb_s1_writedata;                                            // mm_interconnect_1:usb_s1_writedata -> usb:avs_s1_writedata
	wire         mm_interconnect_1_systimer_s1_chipselect;                                      // mm_interconnect_1:systimer_s1_chipselect -> systimer:chipselect
	wire  [15:0] mm_interconnect_1_systimer_s1_readdata;                                        // systimer:readdata -> mm_interconnect_1:systimer_s1_readdata
	wire   [2:0] mm_interconnect_1_systimer_s1_address;                                         // mm_interconnect_1:systimer_s1_address -> systimer:address
	wire         mm_interconnect_1_systimer_s1_write;                                           // mm_interconnect_1:systimer_s1_write -> systimer:write_n
	wire  [15:0] mm_interconnect_1_systimer_s1_writedata;                                       // mm_interconnect_1:systimer_s1_writedata -> systimer:writedata
	wire         mm_interconnect_1_led_s1_chipselect;                                           // mm_interconnect_1:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_1_led_s1_readdata;                                             // led:readdata -> mm_interconnect_1:led_s1_readdata
	wire   [1:0] mm_interconnect_1_led_s1_address;                                              // mm_interconnect_1:led_s1_address -> led:address
	wire         mm_interconnect_1_led_s1_write;                                                // mm_interconnect_1:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_1_led_s1_writedata;                                            // mm_interconnect_1:led_s1_writedata -> led:writedata
	wire         mm_interconnect_1_led_7seg_0_s1_chipselect;                                    // mm_interconnect_1:led_7seg_0_s1_chipselect -> led_7seg_0:chipselect
	wire  [31:0] mm_interconnect_1_led_7seg_0_s1_readdata;                                      // led_7seg_0:readdata -> mm_interconnect_1:led_7seg_0_s1_readdata
	wire   [1:0] mm_interconnect_1_led_7seg_0_s1_address;                                       // mm_interconnect_1:led_7seg_0_s1_address -> led_7seg_0:address
	wire         mm_interconnect_1_led_7seg_0_s1_write;                                         // mm_interconnect_1:led_7seg_0_s1_write -> led_7seg_0:write_n
	wire  [31:0] mm_interconnect_1_led_7seg_0_s1_writedata;                                     // mm_interconnect_1:led_7seg_0_s1_writedata -> led_7seg_0:writedata
	wire         mm_interconnect_1_led_7seg_1_s1_chipselect;                                    // mm_interconnect_1:led_7seg_1_s1_chipselect -> led_7seg_1:chipselect
	wire  [31:0] mm_interconnect_1_led_7seg_1_s1_readdata;                                      // led_7seg_1:readdata -> mm_interconnect_1:led_7seg_1_s1_readdata
	wire   [1:0] mm_interconnect_1_led_7seg_1_s1_address;                                       // mm_interconnect_1:led_7seg_1_s1_address -> led_7seg_1:address
	wire         mm_interconnect_1_led_7seg_1_s1_write;                                         // mm_interconnect_1:led_7seg_1_s1_write -> led_7seg_1:write_n
	wire  [31:0] mm_interconnect_1_led_7seg_1_s1_writedata;                                     // mm_interconnect_1:led_7seg_1_s1_writedata -> led_7seg_1:writedata
	wire         mm_interconnect_1_led_7seg_2_s1_chipselect;                                    // mm_interconnect_1:led_7seg_2_s1_chipselect -> led_7seg_2:chipselect
	wire  [31:0] mm_interconnect_1_led_7seg_2_s1_readdata;                                      // led_7seg_2:readdata -> mm_interconnect_1:led_7seg_2_s1_readdata
	wire   [1:0] mm_interconnect_1_led_7seg_2_s1_address;                                       // mm_interconnect_1:led_7seg_2_s1_address -> led_7seg_2:address
	wire         mm_interconnect_1_led_7seg_2_s1_write;                                         // mm_interconnect_1:led_7seg_2_s1_write -> led_7seg_2:write_n
	wire  [31:0] mm_interconnect_1_led_7seg_2_s1_writedata;                                     // mm_interconnect_1:led_7seg_2_s1_writedata -> led_7seg_2:writedata
	wire         mm_interconnect_1_psw_s1_chipselect;                                           // mm_interconnect_1:psw_s1_chipselect -> psw:chipselect
	wire  [31:0] mm_interconnect_1_psw_s1_readdata;                                             // psw:readdata -> mm_interconnect_1:psw_s1_readdata
	wire   [1:0] mm_interconnect_1_psw_s1_address;                                              // mm_interconnect_1:psw_s1_address -> psw:address
	wire         mm_interconnect_1_psw_s1_write;                                                // mm_interconnect_1:psw_s1_write -> psw:write_n
	wire  [31:0] mm_interconnect_1_psw_s1_writedata;                                            // mm_interconnect_1:psw_s1_writedata -> psw:writedata
	wire  [31:0] mm_interconnect_1_dipsw_s1_readdata;                                           // dipsw:readdata -> mm_interconnect_1:dipsw_s1_readdata
	wire   [1:0] mm_interconnect_1_dipsw_s1_address;                                            // mm_interconnect_1:dipsw_s1_address -> dipsw:address
	wire         mm_interconnect_1_gpio0_s1_chipselect;                                         // mm_interconnect_1:gpio0_s1_chipselect -> gpio0:chipselect
	wire  [31:0] mm_interconnect_1_gpio0_s1_readdata;                                           // gpio0:readdata -> mm_interconnect_1:gpio0_s1_readdata
	wire   [1:0] mm_interconnect_1_gpio0_s1_address;                                            // mm_interconnect_1:gpio0_s1_address -> gpio0:address
	wire         mm_interconnect_1_gpio0_s1_write;                                              // mm_interconnect_1:gpio0_s1_write -> gpio0:write_n
	wire  [31:0] mm_interconnect_1_gpio0_s1_writedata;                                          // mm_interconnect_1:gpio0_s1_writedata -> gpio0:writedata
	wire         mm_interconnect_1_mmcdma_s1_chipselect;                                        // mm_interconnect_1:mmcdma_s1_chipselect -> mmcdma:chipselect
	wire  [31:0] mm_interconnect_1_mmcdma_s1_readdata;                                          // mmcdma:readdata -> mm_interconnect_1:mmcdma_s1_readdata
	wire   [7:0] mm_interconnect_1_mmcdma_s1_address;                                           // mm_interconnect_1:mmcdma_s1_address -> mmcdma:address
	wire         mm_interconnect_1_mmcdma_s1_read;                                              // mm_interconnect_1:mmcdma_s1_read -> mmcdma:read
	wire         mm_interconnect_1_mmcdma_s1_write;                                             // mm_interconnect_1:mmcdma_s1_write -> mmcdma:write
	wire  [31:0] mm_interconnect_1_mmcdma_s1_writedata;                                         // mm_interconnect_1:mmcdma_s1_writedata -> mmcdma:writedata
	wire  [31:0] nios2_fast_irq_irq;                                                            // irq_mapper:sender_irq -> nios2_fast:irq
	wire         irq_mapper_receiver0_irq;                                                      // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                                 // ps2_kb:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                                      // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                                             // mmcdma:irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver2_irq;                                                      // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                                             // epcq:irq -> irq_synchronizer_002:receiver_irq
	wire         irq_mapper_receiver3_irq;                                                      // irq_synchronizer_003:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_003_receiver_irq;                                             // vga:irq_s1 -> irq_synchronizer_003:receiver_irq
	wire         irq_mapper_receiver4_irq;                                                      // irq_synchronizer_004:sender_irq -> irq_mapper:receiver4_irq
	wire   [0:0] irq_synchronizer_004_receiver_irq;                                             // systimer:irq -> irq_synchronizer_004:receiver_irq
	wire         irq_mapper_receiver5_irq;                                                      // irq_synchronizer_005:sender_irq -> irq_mapper:receiver5_irq
	wire   [0:0] irq_synchronizer_005_receiver_irq;                                             // jtag_uart:av_irq -> irq_synchronizer_005:receiver_irq
	wire         irq_mapper_receiver6_irq;                                                      // irq_synchronizer_006:sender_irq -> irq_mapper:receiver6_irq
	wire   [0:0] irq_synchronizer_006_receiver_irq;                                             // psw:irq -> irq_synchronizer_006:receiver_irq
	wire         irq_mapper_receiver7_irq;                                                      // irq_synchronizer_007:sender_irq -> irq_mapper:receiver7_irq
	wire   [0:0] irq_synchronizer_007_receiver_irq;                                             // usb:avs_s1_irq -> irq_synchronizer_007:receiver_irq
	wire         irq_mapper_receiver8_irq;                                                      // irq_synchronizer_008:sender_irq -> irq_mapper:receiver8_irq
	wire   [0:0] irq_synchronizer_008_receiver_irq;                                             // pcm:ins_irq -> irq_synchronizer_008:receiver_irq
	wire         rst_controller_reset_out_reset;                                                // rst_controller:reset_out -> [bootmem:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, irq_synchronizer_005:sender_reset, irq_synchronizer_006:sender_reset, irq_synchronizer_007:sender_reset, irq_synchronizer_008:sender_reset, mm_interconnect_0:nios2_fast_reset_reset_bridge_in_reset_reset, nios2_fast:reset_n, peripherals_bridge:s0_reset, rst_translator:in_reset, sdram:reset_n]
	wire         rst_controller_reset_out_reset_req;                                            // rst_controller:reset_req -> [bootmem:reset_req, nios2_fast:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                            // rst_controller_001:reset_out -> [dipsw:reset_n, epcq:reset_n, gpio0:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, irq_synchronizer_004:receiver_reset, irq_synchronizer_005:receiver_reset, irq_synchronizer_006:receiver_reset, irq_synchronizer_007:receiver_reset, irq_synchronizer_008:receiver_reset, jtag_uart:rst_n, led:reset_n, led_7seg_0:reset_n, led_7seg_1:reset_n, led_7seg_2:reset_n, mm_interconnect_1:peripherals_bridge_m0_reset_reset_bridge_in_reset_reset, mmcdma:reset, pcm:csi_reset, peripherals_bridge:m0_reset, ps2_kb:reset, psw:reset_n, sysid:reset_n, systimer:reset_n, usb:avs_s1_reset, vga:g_reset]
	wire         rst_controller_002_reset_out_reset;                                            // rst_controller_002:reset_out -> mm_interconnect_0:vga_g_reset_reset_bridge_in_reset_reset

	cineraria_core_bootmem bootmem (
		.clk        (core_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_bootmem_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_bootmem_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_bootmem_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_bootmem_s1_write),      //       .write
		.readdata   (mm_interconnect_0_bootmem_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_bootmem_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_bootmem_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),          // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)       //       .reset_req
	);

	cineraria_core_dipsw dipsw (
		.clk      (peri_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_1_dipsw_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_dipsw_s1_readdata), //                    .readdata
		.in_port  (dipsw_export)                         // external_connection.export
	);

	altera_epcq_controller_wrapper #(
		.DEVICE_FAMILY     ("Cyclone V"),
		.ASI_WIDTH         (1),
		.CS_WIDTH          (1),
		.ADDR_WIDTH        (21),
		.ASMI_ADDR_WIDTH   (24),
		.ENABLE_4BYTE_ADDR (0),
		.CHIP_SELS         (1)
	) epcq (
		.clk                  (peri_clk),                                     //       clock_sink.clk
		.reset_n              (~rst_controller_001_reset_out_reset),          //            reset.reset_n
		.avl_csr_read         (mm_interconnect_1_epcq_avl_csr_read),          //          avl_csr.read
		.avl_csr_waitrequest  (mm_interconnect_1_epcq_avl_csr_waitrequest),   //                 .waitrequest
		.avl_csr_write        (mm_interconnect_1_epcq_avl_csr_write),         //                 .write
		.avl_csr_addr         (mm_interconnect_1_epcq_avl_csr_address),       //                 .address
		.avl_csr_wrdata       (mm_interconnect_1_epcq_avl_csr_writedata),     //                 .writedata
		.avl_csr_rddata       (mm_interconnect_1_epcq_avl_csr_readdata),      //                 .readdata
		.avl_csr_rddata_valid (mm_interconnect_1_epcq_avl_csr_readdatavalid), //                 .readdatavalid
		.avl_mem_write        (mm_interconnect_1_epcq_avl_mem_write),         //          avl_mem.write
		.avl_mem_burstcount   (mm_interconnect_1_epcq_avl_mem_burstcount),    //                 .burstcount
		.avl_mem_waitrequest  (mm_interconnect_1_epcq_avl_mem_waitrequest),   //                 .waitrequest
		.avl_mem_read         (mm_interconnect_1_epcq_avl_mem_read),          //                 .read
		.avl_mem_addr         (mm_interconnect_1_epcq_avl_mem_address),       //                 .address
		.avl_mem_wrdata       (mm_interconnect_1_epcq_avl_mem_writedata),     //                 .writedata
		.avl_mem_rddata       (mm_interconnect_1_epcq_avl_mem_readdata),      //                 .readdata
		.avl_mem_rddata_valid (mm_interconnect_1_epcq_avl_mem_readdatavalid), //                 .readdatavalid
		.avl_mem_byteenable   (mm_interconnect_1_epcq_avl_mem_byteenable),    //                 .byteenable
		.irq                  (irq_synchronizer_002_receiver_irq)             // interrupt_sender.irq
	);

	cineraria_core_gpio0 gpio0 (
		.clk        (peri_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address    (mm_interconnect_1_gpio0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_gpio0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_gpio0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_gpio0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_gpio0_s1_readdata),   //                    .readdata
		.bidir_port (gpio0_export)                           // external_connection.export
	);

	cineraria_core_jtag_uart jtag_uart (
		.clk            (peri_clk),                                                  //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_005_receiver_irq)                          //               irq.irq
	);

	cineraria_core_led led (
		.clk        (peri_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                           // external_connection.export
	);

	cineraria_core_led_7seg_0 led_7seg_0 (
		.clk        (peri_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_1_led_7seg_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_7seg_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_7seg_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_7seg_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_7seg_0_s1_readdata),   //                    .readdata
		.out_port   (led7seg_0_export)                            // external_connection.export
	);

	cineraria_core_led_7seg_0 led_7seg_1 (
		.clk        (peri_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_1_led_7seg_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_7seg_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_7seg_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_7seg_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_7seg_1_s1_readdata),   //                    .readdata
		.out_port   (led7seg_1_export)                            // external_connection.export
	);

	cineraria_core_led_7seg_0 led_7seg_2 (
		.clk        (peri_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_1_led_7seg_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_7seg_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_7seg_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_7seg_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_7seg_2_s1_readdata),   //                    .readdata
		.out_port   (led7seg_2_export)                            // external_connection.export
	);

	avalonif_mmcdma #(
		.SYSTEMCLOCKINFO (50000000)
	) mmcdma (
		.clk        (peri_clk),                               //       clock_reset.clk
		.reset      (rst_controller_001_reset_out_reset),     // clock_reset_reset.reset
		.chipselect (mm_interconnect_1_mmcdma_s1_chipselect), //                s1.chipselect
		.address    (mm_interconnect_1_mmcdma_s1_address),    //                  .address
		.read       (mm_interconnect_1_mmcdma_s1_read),       //                  .read
		.readdata   (mm_interconnect_1_mmcdma_s1_readdata),   //                  .readdata
		.write      (mm_interconnect_1_mmcdma_s1_write),      //                  .write
		.writedata  (mm_interconnect_1_mmcdma_s1_writedata),  //                  .writedata
		.MMC_nCS    (sd_nCS),                                 //       conduit_end.export
		.MMC_SCK    (sd_SCK),                                 //                  .export
		.MMC_SDO    (sd_SDO),                                 //                  .export
		.MMC_SDI    (sd_SDI),                                 //                  .export
		.MMC_CD     (sd_CD),                                  //                  .export
		.MMC_WP     (sd_WP),                                  //                  .export
		.irq        (irq_synchronizer_001_receiver_irq)       //  interrupt_sender.irq
	);

	cineraria_core_nios2_fast nios2_fast (
		.clk                                 (core_clk),                                                 //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                          //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                       //                          .reset_req
		.d_address                           (nios2_fast_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_fast_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_fast_data_master_read),                              //                          .read
		.d_readdata                          (nios2_fast_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_fast_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_fast_data_master_write),                             //                          .write
		.d_writedata                         (nios2_fast_data_master_writedata),                         //                          .writedata
		.d_burstcount                        (nios2_fast_data_master_burstcount),                        //                          .burstcount
		.d_readdatavalid                     (nios2_fast_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_fast_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_fast_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_fast_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_fast_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_fast_instruction_master_waitrequest),                //                          .waitrequest
		.i_burstcount                        (nios2_fast_instruction_master_burstcount),                 //                          .burstcount
		.i_readdatavalid                     (nios2_fast_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_fast_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                         //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_fast_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_fast_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_fast_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_fast_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_fast_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_fast_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_fast_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_fast_debug_mem_slave_writedata),   //                          .writedata
		.A_ci_multi_done                     (nios2_fast_custom_instruction_master_done),                // custom_instruction_master.done
		.A_ci_multi_result                   (nios2_fast_custom_instruction_master_multi_result),        //                          .multi_result
		.A_ci_multi_a                        (nios2_fast_custom_instruction_master_multi_a),             //                          .multi_a
		.A_ci_multi_b                        (nios2_fast_custom_instruction_master_multi_b),             //                          .multi_b
		.A_ci_multi_c                        (nios2_fast_custom_instruction_master_multi_c),             //                          .multi_c
		.A_ci_multi_clk_en                   (nios2_fast_custom_instruction_master_clk_en),              //                          .clk_en
		.A_ci_multi_clock                    (nios2_fast_custom_instruction_master_clk),                 //                          .clk
		.A_ci_multi_reset                    (nios2_fast_custom_instruction_master_reset),               //                          .reset
		.A_ci_multi_reset_req                (nios2_fast_custom_instruction_master_reset_req),           //                          .reset_req
		.A_ci_multi_dataa                    (nios2_fast_custom_instruction_master_multi_dataa),         //                          .multi_dataa
		.A_ci_multi_datab                    (nios2_fast_custom_instruction_master_multi_datab),         //                          .multi_datab
		.A_ci_multi_n                        (nios2_fast_custom_instruction_master_multi_n),             //                          .multi_n
		.A_ci_multi_readra                   (nios2_fast_custom_instruction_master_multi_readra),        //                          .multi_readra
		.A_ci_multi_readrb                   (nios2_fast_custom_instruction_master_multi_readrb),        //                          .multi_readrb
		.A_ci_multi_start                    (nios2_fast_custom_instruction_master_start),               //                          .start
		.A_ci_multi_writerc                  (nios2_fast_custom_instruction_master_multi_writerc)        //                          .multi_writerc
	);

	fpoint_wrapper #(
		.useDivider (1)
	) nios_custom_instr_floating_point_0 (
		.clk    (nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_clk),    // s1.clk
		.clk_en (nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //   .clk_en
		.dataa  (nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  //   .dataa
		.datab  (nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //   .datab
		.n      (nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_n),      //   .n
		.reset  (nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //   .reset
		.start  (nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_start),  //   .start
		.done   (nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_done),   //   .done
		.result (nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_result)  //   .result
	);

	pcm_component pcm (
		.csi_clk       (peri_clk),                           //  clock.clk
		.avs_address   (mm_interconnect_1_pcm_s0_address),   //     s0.address
		.avs_read      (mm_interconnect_1_pcm_s0_read),      //       .read
		.avs_readdata  (mm_interconnect_1_pcm_s0_readdata),  //       .readdata
		.avs_write     (mm_interconnect_1_pcm_s0_write),     //       .write
		.avs_writedata (mm_interconnect_1_pcm_s0_writedata), //       .writedata
		.csi_reset     (rst_controller_001_reset_out_reset), //  reset.reset
		.ins_irq       (irq_synchronizer_008_receiver_irq),  //    irs.irq
		.coe_aud_clk   (pcm_clk),                            // export.clk
		.coe_aud_mute  (pcm_mute),                           //       .mute
		.coe_aud_l     (pcm_aud_l),                          //       .aud_l
		.coe_aud_r     (pcm_aud_r)                           //       .aud_r
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (24),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) peripherals_bridge (
		.m0_clk           (peri_clk),                                              //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                    // m0_reset.reset
		.s0_clk           (core_clk),                                              //   s0_clk.clk
		.s0_reset         (rst_controller_reset_out_reset),                        // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_peripherals_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_peripherals_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_peripherals_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_peripherals_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_peripherals_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_peripherals_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_peripherals_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_peripherals_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_peripherals_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_peripherals_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (peripherals_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (peripherals_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (peripherals_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (peripherals_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (peripherals_bridge_m0_writedata),                       //         .writedata
		.m0_address       (peripherals_bridge_m0_address),                         //         .address
		.m0_write         (peripherals_bridge_m0_write),                           //         .write
		.m0_read          (peripherals_bridge_m0_read),                            //         .read
		.m0_byteenable    (peripherals_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (peripherals_bridge_m0_debugaccess)                      //         .debugaccess
	);

	pixelsimd pixelsimd (
		.dataa  (nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_dataa),  // nios_custom_instruction_slave_0.dataa
		.datab  (nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_datab),  //                                .datab
		.result (nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_result), //                                .result
		.clk    (nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_clk),    //                                .clk
		.clk_en (nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_clk_en), //                                .clk_en
		.reset  (nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_reset),  //                                .reset
		.start  (nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_start),  //                                .start
		.done   (nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_done),   //                                .done
		.n      (nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_n)       //                                .n
	);

	cineraria_core_ps2_kb ps2_kb (
		.clk         (peri_clk),                                              //                clk.clk
		.reset       (rst_controller_001_reset_out_reset),                    //              reset.reset
		.address     (mm_interconnect_1_ps2_kb_avalon_ps2_slave_address),     //   avalon_ps2_slave.address
		.chipselect  (mm_interconnect_1_ps2_kb_avalon_ps2_slave_chipselect),  //                   .chipselect
		.byteenable  (mm_interconnect_1_ps2_kb_avalon_ps2_slave_byteenable),  //                   .byteenable
		.read        (mm_interconnect_1_ps2_kb_avalon_ps2_slave_read),        //                   .read
		.write       (mm_interconnect_1_ps2_kb_avalon_ps2_slave_write),       //                   .write
		.writedata   (mm_interconnect_1_ps2_kb_avalon_ps2_slave_writedata),   //                   .writedata
		.readdata    (mm_interconnect_1_ps2_kb_avalon_ps2_slave_readdata),    //                   .readdata
		.waitrequest (mm_interconnect_1_ps2_kb_avalon_ps2_slave_waitrequest), //                   .waitrequest
		.irq         (irq_synchronizer_receiver_irq),                         //          interrupt.irq
		.PS2_CLK     (ps2_kb_CLK),                                            // external_interface.export
		.PS2_DAT     (ps2_kb_DAT)                                             //                   .export
	);

	cineraria_core_psw psw (
		.clk        (peri_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_psw_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_psw_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_psw_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_psw_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_psw_s1_readdata),   //                    .readdata
		.in_port    (psw_export),                          // external_connection.export
		.irq        (irq_synchronizer_006_receiver_irq)    //                 irq.irq
	);

	cineraria_core_sdram sdram (
		.clk            (core_clk),                                 //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdr_addr),                                 //  wire.export
		.zs_ba          (sdr_ba),                                   //      .export
		.zs_cas_n       (sdr_cas_n),                                //      .export
		.zs_cke         (sdr_cke),                                  //      .export
		.zs_cs_n        (sdr_cs_n),                                 //      .export
		.zs_dq          (sdr_dq),                                   //      .export
		.zs_dqm         (sdr_dqm),                                  //      .export
		.zs_ras_n       (sdr_ras_n),                                //      .export
		.zs_we_n        (sdr_we_n)                                  //      .export
	);

	cineraria_core_sysid sysid (
		.clock    (peri_clk),                                       //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	cineraria_core_systimer systimer (
		.clk        (peri_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.address    (mm_interconnect_1_systimer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_systimer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_systimer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_systimer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_systimer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_004_receiver_irq)         //   irq.irq
	);

	usbhost_component #(
		.HOST_FIFO_DEPTH      (64),
		.HOST_FIFO_ADDR_WIDTH (6)
	) usb (
		.avs_s1_chipselect  (mm_interconnect_1_usb_s1_chipselect),  //       s1.chipselect
		.avs_s1_address     (mm_interconnect_1_usb_s1_address),     //         .address
		.avs_s1_read        (mm_interconnect_1_usb_s1_read),        //         .read
		.avs_s1_readdata    (mm_interconnect_1_usb_s1_readdata),    //         .readdata
		.avs_s1_write       (mm_interconnect_1_usb_s1_write),       //         .write
		.avs_s1_writedata   (mm_interconnect_1_usb_s1_writedata),   //         .writedata
		.avs_s1_waitrequest (mm_interconnect_1_usb_s1_waitrequest), //         .waitrequest
		.avs_s1_irq         (irq_synchronizer_007_receiver_irq),    //   irq_s1.irq
		.test_dataouttick   (usb_test_dataouttick),                 //  usbport.export
		.test_dataintick    (usb_test_dataintick),                  //         .export
		.usbclk_48mhz       (usb_usbclk_48mhz),                     //         .export
		.usb_dp             (usb_usb_dp),                           //         .export
		.usb_dm             (usb_usb_dm),                           //         .export
		.usb_oe_n           (usb_usb_oe_n),                         //         .export
		.usb_fullspeed      (usb_usb_fullspeed),                    //         .export
		.avs_s1_clk         (peri_clk),                             // clock_s1.clk
		.avs_s1_reset       (rst_controller_001_reset_out_reset)    // reset_s1.reset
	);

	vga_component #(
		.LINEOFFSETBYTES (2048),
		.H_TOTAL         (800),
		.H_SYNC          (96),
		.H_BACKP         (48),
		.H_ACTIVE        (640),
		.V_TOTAL         (525),
		.V_SYNC          (2),
		.V_BACKP         (33),
		.V_ACTIVE        (480)
	) vga (
		.video_clk            (vga_clk),                            //     ext.export
		.video_rout           (vga_rout),                           //        .export
		.video_gout           (vga_gout),                           //        .export
		.video_bout           (vga_bout),                           //        .export
		.video_hsync_n        (vga_hsync_n),                        //        .export
		.video_vsync_n        (vga_vsync_n),                        //        .export
		.video_enable         (vga_enable),                         //        .export
		.avm_m1_address       (vga_m1_address),                     //      m1.address
		.avm_m1_waitrequest   (vga_m1_waitrequest),                 //        .waitrequest
		.avm_m1_burstcount    (vga_m1_burstcount),                  //        .burstcount
		.avm_m1_read          (vga_m1_read),                        //        .read
		.avm_m1_readdata      (vga_m1_readdata),                    //        .readdata
		.avm_m1_readdatavalid (vga_m1_readdatavalid),               //        .readdatavalid
		.avs_s1_address       (mm_interconnect_1_vga_s1_address),   //      s1.address
		.avs_s1_read          (mm_interconnect_1_vga_s1_read),      //        .read
		.avs_s1_readdata      (mm_interconnect_1_vga_s1_readdata),  //        .readdata
		.avs_s1_write         (mm_interconnect_1_vga_s1_write),     //        .write
		.avs_s1_writedata     (mm_interconnect_1_vga_s1_writedata), //        .writedata
		.irq_s1               (irq_synchronizer_003_receiver_irq),  //     irq.irq
		.s1_clk               (peri_clk),                           //   s_clk.clk
		.m1_clk               (core_clk),                           //   m_clk.clk
		.g_reset              (rst_controller_001_reset_out_reset)  // g_reset.reset
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) nios2_fast_custom_instruction_master_translator (
		.ci_slave_result           (),                                                                          //        ci_slave.result
		.ci_slave_multi_clk        (nios2_fast_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios2_fast_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios2_fast_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios2_fast_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios2_fast_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios2_fast_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (nios2_fast_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (nios2_fast_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (nios2_fast_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (nios2_fast_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (nios2_fast_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (nios2_fast_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (nios2_fast_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (nios2_fast_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (nios2_fast_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (nios2_fast_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_result     (),                                                                          //  comb_ci_master.result
		.multi_ci_master_clk       (nios2_fast_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios2_fast_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios2_fast_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios2_fast_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios2_fast_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios2_fast_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios2_fast_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios2_fast_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios2_fast_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios2_fast_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios2_fast_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios2_fast_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios2_fast_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios2_fast_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios2_fast_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios2_fast_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_dataa            (32'b00000000000000000000000000000000),                                      //     (terminated)
		.ci_slave_datab            (32'b00000000000000000000000000000000),                                      //     (terminated)
		.ci_slave_n                (8'b00000000),                                                               //     (terminated)
		.ci_slave_readra           (1'b0),                                                                      //     (terminated)
		.ci_slave_readrb           (1'b0),                                                                      //     (terminated)
		.ci_slave_writerc          (1'b0),                                                                      //     (terminated)
		.ci_slave_a                (5'b00000),                                                                  //     (terminated)
		.ci_slave_b                (5'b00000),                                                                  //     (terminated)
		.ci_slave_c                (5'b00000),                                                                  //     (terminated)
		.ci_slave_ipending         (32'b00000000000000000000000000000000),                                      //     (terminated)
		.ci_slave_estatus          (1'b0),                                                                      //     (terminated)
		.comb_ci_master_dataa      (),                                                                          //     (terminated)
		.comb_ci_master_datab      (),                                                                          //     (terminated)
		.comb_ci_master_n          (),                                                                          //     (terminated)
		.comb_ci_master_readra     (),                                                                          //     (terminated)
		.comb_ci_master_readrb     (),                                                                          //     (terminated)
		.comb_ci_master_writerc    (),                                                                          //     (terminated)
		.comb_ci_master_a          (),                                                                          //     (terminated)
		.comb_ci_master_b          (),                                                                          //     (terminated)
		.comb_ci_master_c          (),                                                                          //     (terminated)
		.comb_ci_master_ipending   (),                                                                          //     (terminated)
		.comb_ci_master_estatus    ()                                                                           //     (terminated)
	);

	cineraria_core_nios2_fast_custom_instruction_master_multi_xconnect nios2_fast_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios2_fast_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios2_fast_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios2_fast_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios2_fast_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios2_fast_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios2_fast_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios2_fast_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios2_fast_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios2_fast_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios2_fast_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                          //           .ipending
		.ci_slave_estatus     (),                                                                          //           .estatus
		.ci_slave_clk         (nios2_fast_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios2_fast_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios2_fast_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios2_fast_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios2_fast_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios2_fast_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_done),       //           .done
		.ci_master1_dataa     (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_dataa),      // ci_master1.dataa
		.ci_master1_datab     (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_datab),      //           .datab
		.ci_master1_result    (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_result),     //           .result
		.ci_master1_n         (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_n),          //           .n
		.ci_master1_readra    (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_readra),     //           .readra
		.ci_master1_readrb    (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_readrb),     //           .readrb
		.ci_master1_writerc   (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_writerc),    //           .writerc
		.ci_master1_a         (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_a),          //           .a
		.ci_master1_b         (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_b),          //           .b
		.ci_master1_c         (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_c),          //           .c
		.ci_master1_ipending  (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_ipending),   //           .ipending
		.ci_master1_estatus   (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_estatus),    //           .estatus
		.ci_master1_clk       (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_clk),        //           .clk
		.ci_master1_reset     (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_reset),      //           .reset
		.ci_master1_clken     (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_clk_en),     //           .clk_en
		.ci_master1_reset_req (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_reset_req),  //           .reset_req
		.ci_master1_start     (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_start),      //           .start
		.ci_master1_done      (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (2),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) nios2_fast_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_n),      //          .n
		.ci_master_clk       (nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_readra    (),                                                                              // (terminated)
		.ci_master_readrb    (),                                                                              // (terminated)
		.ci_master_writerc   (),                                                                              // (terminated)
		.ci_master_a         (),                                                                              // (terminated)
		.ci_master_b         (),                                                                              // (terminated)
		.ci_master_c         (),                                                                              // (terminated)
		.ci_master_ipending  (),                                                                              // (terminated)
		.ci_master_estatus   (),                                                                              // (terminated)
		.ci_master_reset_req ()                                                                               // (terminated)
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios2_fast_custom_instruction_master_multi_slave_translator1 (
		.ci_slave_dataa      (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_datab),          //          .datab
		.ci_slave_result     (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_result),         //          .result
		.ci_slave_n          (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_n),              //          .n
		.ci_slave_readra     (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_readra),         //          .readra
		.ci_slave_readrb     (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_writerc),        //          .writerc
		.ci_slave_a          (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_a),              //          .a
		.ci_slave_b          (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_b),              //          .b
		.ci_slave_c          (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_c),              //          .c
		.ci_slave_ipending   (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_estatus),        //          .estatus
		.ci_slave_clk        (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_clk),            //          .clk
		.ci_slave_clken      (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_reset),          //          .reset
		.ci_slave_start      (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_start),          //          .start
		.ci_slave_done       (nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_done),           //          .done
		.ci_master_dataa     (nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_result), //          .result
		.ci_master_n         (nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_n),      //          .n
		.ci_master_clk       (nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_reset),  //          .reset
		.ci_master_start     (nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_start),  //          .start
		.ci_master_done      (nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_done),   //          .done
		.ci_master_readra    (),                                                                              // (terminated)
		.ci_master_readrb    (),                                                                              // (terminated)
		.ci_master_writerc   (),                                                                              // (terminated)
		.ci_master_a         (),                                                                              // (terminated)
		.ci_master_b         (),                                                                              // (terminated)
		.ci_master_c         (),                                                                              // (terminated)
		.ci_master_ipending  (),                                                                              // (terminated)
		.ci_master_estatus   (),                                                                              // (terminated)
		.ci_master_reset_req ()                                                                               // (terminated)
	);

	cineraria_core_mm_interconnect_0 mm_interconnect_0 (
		.clk_core_clk_clk                             (core_clk),                                                 //                           clk_core_clk.clk
		.nios2_fast_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                           // nios2_fast_reset_reset_bridge_in_reset.reset
		.vga_g_reset_reset_bridge_in_reset_reset      (rst_controller_002_reset_out_reset),                       //      vga_g_reset_reset_bridge_in_reset.reset
		.nios2_fast_data_master_address               (nios2_fast_data_master_address),                           //                 nios2_fast_data_master.address
		.nios2_fast_data_master_waitrequest           (nios2_fast_data_master_waitrequest),                       //                                       .waitrequest
		.nios2_fast_data_master_burstcount            (nios2_fast_data_master_burstcount),                        //                                       .burstcount
		.nios2_fast_data_master_byteenable            (nios2_fast_data_master_byteenable),                        //                                       .byteenable
		.nios2_fast_data_master_read                  (nios2_fast_data_master_read),                              //                                       .read
		.nios2_fast_data_master_readdata              (nios2_fast_data_master_readdata),                          //                                       .readdata
		.nios2_fast_data_master_readdatavalid         (nios2_fast_data_master_readdatavalid),                     //                                       .readdatavalid
		.nios2_fast_data_master_write                 (nios2_fast_data_master_write),                             //                                       .write
		.nios2_fast_data_master_writedata             (nios2_fast_data_master_writedata),                         //                                       .writedata
		.nios2_fast_data_master_debugaccess           (nios2_fast_data_master_debugaccess),                       //                                       .debugaccess
		.nios2_fast_instruction_master_address        (nios2_fast_instruction_master_address),                    //          nios2_fast_instruction_master.address
		.nios2_fast_instruction_master_waitrequest    (nios2_fast_instruction_master_waitrequest),                //                                       .waitrequest
		.nios2_fast_instruction_master_burstcount     (nios2_fast_instruction_master_burstcount),                 //                                       .burstcount
		.nios2_fast_instruction_master_read           (nios2_fast_instruction_master_read),                       //                                       .read
		.nios2_fast_instruction_master_readdata       (nios2_fast_instruction_master_readdata),                   //                                       .readdata
		.nios2_fast_instruction_master_readdatavalid  (nios2_fast_instruction_master_readdatavalid),              //                                       .readdatavalid
		.vga_m1_address                               (vga_m1_address),                                           //                                 vga_m1.address
		.vga_m1_waitrequest                           (vga_m1_waitrequest),                                       //                                       .waitrequest
		.vga_m1_burstcount                            (vga_m1_burstcount),                                        //                                       .burstcount
		.vga_m1_read                                  (vga_m1_read),                                              //                                       .read
		.vga_m1_readdata                              (vga_m1_readdata),                                          //                                       .readdata
		.vga_m1_readdatavalid                         (vga_m1_readdatavalid),                                     //                                       .readdatavalid
		.bootmem_s1_address                           (mm_interconnect_0_bootmem_s1_address),                     //                             bootmem_s1.address
		.bootmem_s1_write                             (mm_interconnect_0_bootmem_s1_write),                       //                                       .write
		.bootmem_s1_readdata                          (mm_interconnect_0_bootmem_s1_readdata),                    //                                       .readdata
		.bootmem_s1_writedata                         (mm_interconnect_0_bootmem_s1_writedata),                   //                                       .writedata
		.bootmem_s1_byteenable                        (mm_interconnect_0_bootmem_s1_byteenable),                  //                                       .byteenable
		.bootmem_s1_chipselect                        (mm_interconnect_0_bootmem_s1_chipselect),                  //                                       .chipselect
		.bootmem_s1_clken                             (mm_interconnect_0_bootmem_s1_clken),                       //                                       .clken
		.nios2_fast_debug_mem_slave_address           (mm_interconnect_0_nios2_fast_debug_mem_slave_address),     //             nios2_fast_debug_mem_slave.address
		.nios2_fast_debug_mem_slave_write             (mm_interconnect_0_nios2_fast_debug_mem_slave_write),       //                                       .write
		.nios2_fast_debug_mem_slave_read              (mm_interconnect_0_nios2_fast_debug_mem_slave_read),        //                                       .read
		.nios2_fast_debug_mem_slave_readdata          (mm_interconnect_0_nios2_fast_debug_mem_slave_readdata),    //                                       .readdata
		.nios2_fast_debug_mem_slave_writedata         (mm_interconnect_0_nios2_fast_debug_mem_slave_writedata),   //                                       .writedata
		.nios2_fast_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_fast_debug_mem_slave_byteenable),  //                                       .byteenable
		.nios2_fast_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_fast_debug_mem_slave_waitrequest), //                                       .waitrequest
		.nios2_fast_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_fast_debug_mem_slave_debugaccess), //                                       .debugaccess
		.peripherals_bridge_s0_address                (mm_interconnect_0_peripherals_bridge_s0_address),          //                  peripherals_bridge_s0.address
		.peripherals_bridge_s0_write                  (mm_interconnect_0_peripherals_bridge_s0_write),            //                                       .write
		.peripherals_bridge_s0_read                   (mm_interconnect_0_peripherals_bridge_s0_read),             //                                       .read
		.peripherals_bridge_s0_readdata               (mm_interconnect_0_peripherals_bridge_s0_readdata),         //                                       .readdata
		.peripherals_bridge_s0_writedata              (mm_interconnect_0_peripherals_bridge_s0_writedata),        //                                       .writedata
		.peripherals_bridge_s0_burstcount             (mm_interconnect_0_peripherals_bridge_s0_burstcount),       //                                       .burstcount
		.peripherals_bridge_s0_byteenable             (mm_interconnect_0_peripherals_bridge_s0_byteenable),       //                                       .byteenable
		.peripherals_bridge_s0_readdatavalid          (mm_interconnect_0_peripherals_bridge_s0_readdatavalid),    //                                       .readdatavalid
		.peripherals_bridge_s0_waitrequest            (mm_interconnect_0_peripherals_bridge_s0_waitrequest),      //                                       .waitrequest
		.peripherals_bridge_s0_debugaccess            (mm_interconnect_0_peripherals_bridge_s0_debugaccess),      //                                       .debugaccess
		.sdram_s1_address                             (mm_interconnect_0_sdram_s1_address),                       //                               sdram_s1.address
		.sdram_s1_write                               (mm_interconnect_0_sdram_s1_write),                         //                                       .write
		.sdram_s1_read                                (mm_interconnect_0_sdram_s1_read),                          //                                       .read
		.sdram_s1_readdata                            (mm_interconnect_0_sdram_s1_readdata),                      //                                       .readdata
		.sdram_s1_writedata                           (mm_interconnect_0_sdram_s1_writedata),                     //                                       .writedata
		.sdram_s1_byteenable                          (mm_interconnect_0_sdram_s1_byteenable),                    //                                       .byteenable
		.sdram_s1_readdatavalid                       (mm_interconnect_0_sdram_s1_readdatavalid),                 //                                       .readdatavalid
		.sdram_s1_waitrequest                         (mm_interconnect_0_sdram_s1_waitrequest),                   //                                       .waitrequest
		.sdram_s1_chipselect                          (mm_interconnect_0_sdram_s1_chipselect)                     //                                       .chipselect
	);

	cineraria_core_mm_interconnect_1 mm_interconnect_1 (
		.clk_peri_clk_clk                                        (peri_clk),                                                  //                                      clk_peri_clk.clk
		.peripherals_bridge_m0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                        // peripherals_bridge_m0_reset_reset_bridge_in_reset.reset
		.peripherals_bridge_m0_address                           (peripherals_bridge_m0_address),                             //                             peripherals_bridge_m0.address
		.peripherals_bridge_m0_waitrequest                       (peripherals_bridge_m0_waitrequest),                         //                                                  .waitrequest
		.peripherals_bridge_m0_burstcount                        (peripherals_bridge_m0_burstcount),                          //                                                  .burstcount
		.peripherals_bridge_m0_byteenable                        (peripherals_bridge_m0_byteenable),                          //                                                  .byteenable
		.peripherals_bridge_m0_read                              (peripherals_bridge_m0_read),                                //                                                  .read
		.peripherals_bridge_m0_readdata                          (peripherals_bridge_m0_readdata),                            //                                                  .readdata
		.peripherals_bridge_m0_readdatavalid                     (peripherals_bridge_m0_readdatavalid),                       //                                                  .readdatavalid
		.peripherals_bridge_m0_write                             (peripherals_bridge_m0_write),                               //                                                  .write
		.peripherals_bridge_m0_writedata                         (peripherals_bridge_m0_writedata),                           //                                                  .writedata
		.peripherals_bridge_m0_debugaccess                       (peripherals_bridge_m0_debugaccess),                         //                                                  .debugaccess
		.dipsw_s1_address                                        (mm_interconnect_1_dipsw_s1_address),                        //                                          dipsw_s1.address
		.dipsw_s1_readdata                                       (mm_interconnect_1_dipsw_s1_readdata),                       //                                                  .readdata
		.epcq_avl_csr_address                                    (mm_interconnect_1_epcq_avl_csr_address),                    //                                      epcq_avl_csr.address
		.epcq_avl_csr_write                                      (mm_interconnect_1_epcq_avl_csr_write),                      //                                                  .write
		.epcq_avl_csr_read                                       (mm_interconnect_1_epcq_avl_csr_read),                       //                                                  .read
		.epcq_avl_csr_readdata                                   (mm_interconnect_1_epcq_avl_csr_readdata),                   //                                                  .readdata
		.epcq_avl_csr_writedata                                  (mm_interconnect_1_epcq_avl_csr_writedata),                  //                                                  .writedata
		.epcq_avl_csr_readdatavalid                              (mm_interconnect_1_epcq_avl_csr_readdatavalid),              //                                                  .readdatavalid
		.epcq_avl_csr_waitrequest                                (mm_interconnect_1_epcq_avl_csr_waitrequest),                //                                                  .waitrequest
		.epcq_avl_mem_address                                    (mm_interconnect_1_epcq_avl_mem_address),                    //                                      epcq_avl_mem.address
		.epcq_avl_mem_write                                      (mm_interconnect_1_epcq_avl_mem_write),                      //                                                  .write
		.epcq_avl_mem_read                                       (mm_interconnect_1_epcq_avl_mem_read),                       //                                                  .read
		.epcq_avl_mem_readdata                                   (mm_interconnect_1_epcq_avl_mem_readdata),                   //                                                  .readdata
		.epcq_avl_mem_writedata                                  (mm_interconnect_1_epcq_avl_mem_writedata),                  //                                                  .writedata
		.epcq_avl_mem_burstcount                                 (mm_interconnect_1_epcq_avl_mem_burstcount),                 //                                                  .burstcount
		.epcq_avl_mem_byteenable                                 (mm_interconnect_1_epcq_avl_mem_byteenable),                 //                                                  .byteenable
		.epcq_avl_mem_readdatavalid                              (mm_interconnect_1_epcq_avl_mem_readdatavalid),              //                                                  .readdatavalid
		.epcq_avl_mem_waitrequest                                (mm_interconnect_1_epcq_avl_mem_waitrequest),                //                                                  .waitrequest
		.gpio0_s1_address                                        (mm_interconnect_1_gpio0_s1_address),                        //                                          gpio0_s1.address
		.gpio0_s1_write                                          (mm_interconnect_1_gpio0_s1_write),                          //                                                  .write
		.gpio0_s1_readdata                                       (mm_interconnect_1_gpio0_s1_readdata),                       //                                                  .readdata
		.gpio0_s1_writedata                                      (mm_interconnect_1_gpio0_s1_writedata),                      //                                                  .writedata
		.gpio0_s1_chipselect                                     (mm_interconnect_1_gpio0_s1_chipselect),                     //                                                  .chipselect
		.jtag_uart_avalon_jtag_slave_address                     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                       jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                       (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),       //                                                  .write
		.jtag_uart_avalon_jtag_slave_read                        (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),        //                                                  .read
		.jtag_uart_avalon_jtag_slave_readdata                    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                                                  .readdata
		.jtag_uart_avalon_jtag_slave_writedata                   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                                                  .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                 (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                                                  .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  //                                                  .chipselect
		.led_s1_address                                          (mm_interconnect_1_led_s1_address),                          //                                            led_s1.address
		.led_s1_write                                            (mm_interconnect_1_led_s1_write),                            //                                                  .write
		.led_s1_readdata                                         (mm_interconnect_1_led_s1_readdata),                         //                                                  .readdata
		.led_s1_writedata                                        (mm_interconnect_1_led_s1_writedata),                        //                                                  .writedata
		.led_s1_chipselect                                       (mm_interconnect_1_led_s1_chipselect),                       //                                                  .chipselect
		.led_7seg_0_s1_address                                   (mm_interconnect_1_led_7seg_0_s1_address),                   //                                     led_7seg_0_s1.address
		.led_7seg_0_s1_write                                     (mm_interconnect_1_led_7seg_0_s1_write),                     //                                                  .write
		.led_7seg_0_s1_readdata                                  (mm_interconnect_1_led_7seg_0_s1_readdata),                  //                                                  .readdata
		.led_7seg_0_s1_writedata                                 (mm_interconnect_1_led_7seg_0_s1_writedata),                 //                                                  .writedata
		.led_7seg_0_s1_chipselect                                (mm_interconnect_1_led_7seg_0_s1_chipselect),                //                                                  .chipselect
		.led_7seg_1_s1_address                                   (mm_interconnect_1_led_7seg_1_s1_address),                   //                                     led_7seg_1_s1.address
		.led_7seg_1_s1_write                                     (mm_interconnect_1_led_7seg_1_s1_write),                     //                                                  .write
		.led_7seg_1_s1_readdata                                  (mm_interconnect_1_led_7seg_1_s1_readdata),                  //                                                  .readdata
		.led_7seg_1_s1_writedata                                 (mm_interconnect_1_led_7seg_1_s1_writedata),                 //                                                  .writedata
		.led_7seg_1_s1_chipselect                                (mm_interconnect_1_led_7seg_1_s1_chipselect),                //                                                  .chipselect
		.led_7seg_2_s1_address                                   (mm_interconnect_1_led_7seg_2_s1_address),                   //                                     led_7seg_2_s1.address
		.led_7seg_2_s1_write                                     (mm_interconnect_1_led_7seg_2_s1_write),                     //                                                  .write
		.led_7seg_2_s1_readdata                                  (mm_interconnect_1_led_7seg_2_s1_readdata),                  //                                                  .readdata
		.led_7seg_2_s1_writedata                                 (mm_interconnect_1_led_7seg_2_s1_writedata),                 //                                                  .writedata
		.led_7seg_2_s1_chipselect                                (mm_interconnect_1_led_7seg_2_s1_chipselect),                //                                                  .chipselect
		.mmcdma_s1_address                                       (mm_interconnect_1_mmcdma_s1_address),                       //                                         mmcdma_s1.address
		.mmcdma_s1_write                                         (mm_interconnect_1_mmcdma_s1_write),                         //                                                  .write
		.mmcdma_s1_read                                          (mm_interconnect_1_mmcdma_s1_read),                          //                                                  .read
		.mmcdma_s1_readdata                                      (mm_interconnect_1_mmcdma_s1_readdata),                      //                                                  .readdata
		.mmcdma_s1_writedata                                     (mm_interconnect_1_mmcdma_s1_writedata),                     //                                                  .writedata
		.mmcdma_s1_chipselect                                    (mm_interconnect_1_mmcdma_s1_chipselect),                    //                                                  .chipselect
		.pcm_s0_address                                          (mm_interconnect_1_pcm_s0_address),                          //                                            pcm_s0.address
		.pcm_s0_write                                            (mm_interconnect_1_pcm_s0_write),                            //                                                  .write
		.pcm_s0_read                                             (mm_interconnect_1_pcm_s0_read),                             //                                                  .read
		.pcm_s0_readdata                                         (mm_interconnect_1_pcm_s0_readdata),                         //                                                  .readdata
		.pcm_s0_writedata                                        (mm_interconnect_1_pcm_s0_writedata),                        //                                                  .writedata
		.ps2_kb_avalon_ps2_slave_address                         (mm_interconnect_1_ps2_kb_avalon_ps2_slave_address),         //                           ps2_kb_avalon_ps2_slave.address
		.ps2_kb_avalon_ps2_slave_write                           (mm_interconnect_1_ps2_kb_avalon_ps2_slave_write),           //                                                  .write
		.ps2_kb_avalon_ps2_slave_read                            (mm_interconnect_1_ps2_kb_avalon_ps2_slave_read),            //                                                  .read
		.ps2_kb_avalon_ps2_slave_readdata                        (mm_interconnect_1_ps2_kb_avalon_ps2_slave_readdata),        //                                                  .readdata
		.ps2_kb_avalon_ps2_slave_writedata                       (mm_interconnect_1_ps2_kb_avalon_ps2_slave_writedata),       //                                                  .writedata
		.ps2_kb_avalon_ps2_slave_byteenable                      (mm_interconnect_1_ps2_kb_avalon_ps2_slave_byteenable),      //                                                  .byteenable
		.ps2_kb_avalon_ps2_slave_waitrequest                     (mm_interconnect_1_ps2_kb_avalon_ps2_slave_waitrequest),     //                                                  .waitrequest
		.ps2_kb_avalon_ps2_slave_chipselect                      (mm_interconnect_1_ps2_kb_avalon_ps2_slave_chipselect),      //                                                  .chipselect
		.psw_s1_address                                          (mm_interconnect_1_psw_s1_address),                          //                                            psw_s1.address
		.psw_s1_write                                            (mm_interconnect_1_psw_s1_write),                            //                                                  .write
		.psw_s1_readdata                                         (mm_interconnect_1_psw_s1_readdata),                         //                                                  .readdata
		.psw_s1_writedata                                        (mm_interconnect_1_psw_s1_writedata),                        //                                                  .writedata
		.psw_s1_chipselect                                       (mm_interconnect_1_psw_s1_chipselect),                       //                                                  .chipselect
		.sysid_control_slave_address                             (mm_interconnect_1_sysid_control_slave_address),             //                               sysid_control_slave.address
		.sysid_control_slave_readdata                            (mm_interconnect_1_sysid_control_slave_readdata),            //                                                  .readdata
		.systimer_s1_address                                     (mm_interconnect_1_systimer_s1_address),                     //                                       systimer_s1.address
		.systimer_s1_write                                       (mm_interconnect_1_systimer_s1_write),                       //                                                  .write
		.systimer_s1_readdata                                    (mm_interconnect_1_systimer_s1_readdata),                    //                                                  .readdata
		.systimer_s1_writedata                                   (mm_interconnect_1_systimer_s1_writedata),                   //                                                  .writedata
		.systimer_s1_chipselect                                  (mm_interconnect_1_systimer_s1_chipselect),                  //                                                  .chipselect
		.usb_s1_address                                          (mm_interconnect_1_usb_s1_address),                          //                                            usb_s1.address
		.usb_s1_write                                            (mm_interconnect_1_usb_s1_write),                            //                                                  .write
		.usb_s1_read                                             (mm_interconnect_1_usb_s1_read),                             //                                                  .read
		.usb_s1_readdata                                         (mm_interconnect_1_usb_s1_readdata),                         //                                                  .readdata
		.usb_s1_writedata                                        (mm_interconnect_1_usb_s1_writedata),                        //                                                  .writedata
		.usb_s1_waitrequest                                      (mm_interconnect_1_usb_s1_waitrequest),                      //                                                  .waitrequest
		.usb_s1_chipselect                                       (mm_interconnect_1_usb_s1_chipselect),                       //                                                  .chipselect
		.vga_s1_address                                          (mm_interconnect_1_vga_s1_address),                          //                                            vga_s1.address
		.vga_s1_write                                            (mm_interconnect_1_vga_s1_write),                            //                                                  .write
		.vga_s1_read                                             (mm_interconnect_1_vga_s1_read),                             //                                                  .read
		.vga_s1_readdata                                         (mm_interconnect_1_vga_s1_readdata),                         //                                                  .readdata
		.vga_s1_writedata                                        (mm_interconnect_1_vga_s1_writedata)                         //                                                  .writedata
	);

	cineraria_core_irq_mapper irq_mapper (
		.clk           (core_clk),                       //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),       // receiver7.irq
		.receiver8_irq (irq_mapper_receiver8_irq),       // receiver8.irq
		.sender_irq    (nios2_fast_irq_irq)              //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (peri_clk),                           //       receiver_clk.clk
		.sender_clk     (core_clk),                           //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (peri_clk),                           //       receiver_clk.clk
		.sender_clk     (core_clk),                           //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (peri_clk),                           //       receiver_clk.clk
		.sender_clk     (core_clk),                           //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (peri_clk),                           //       receiver_clk.clk
		.sender_clk     (core_clk),                           //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_004 (
		.receiver_clk   (peri_clk),                           //       receiver_clk.clk
		.sender_clk     (core_clk),                           //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_004_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_005 (
		.receiver_clk   (peri_clk),                           //       receiver_clk.clk
		.sender_clk     (core_clk),                           //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_005_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver5_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_006 (
		.receiver_clk   (peri_clk),                           //       receiver_clk.clk
		.sender_clk     (core_clk),                           //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_006_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver6_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_007 (
		.receiver_clk   (peri_clk),                           //       receiver_clk.clk
		.sender_clk     (core_clk),                           //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_007_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver7_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_008 (
		.receiver_clk   (peri_clk),                           //       receiver_clk.clk
		.sender_clk     (core_clk),                           //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_008_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver8_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (core_clk),                           //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (peri_clk),                           //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (core_clk),                           //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
